
module BUF(
    input I,
    output O
    );
    assign O=I;
endmodule